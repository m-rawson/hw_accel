package accel_core_pkg;

  // core mem map definition
  
  // memory partitions
  localparam int MMAP_PREPROC_START_ADDR  = 'd0;
  localparam int MMAP_PREPROC_END_ADDR    = 'd1;
  localparam int MMAP_POSTPROC_START_ADDR = 'd2;
  localparam int MMAP_POSTPROC_END_ADDR   = 'd3;
  localparam int MMAP_START_PROC_TRIG     = 'd4;
  
  
  
endpackage 