// core mem

module core_mem #(
)(
  Axi.Slave  mem_bus,
  Axi.Master preproc_data,
  Axi.Slave  postproc_data
);

endmodule