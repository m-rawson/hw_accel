// HW Accelerator wrapper

module hw_accel #(
)(
  input wire    clk,
  input wire    rst,
  Axis.Slave  data_i,
  Axis.Master data_o,
  AXi.Slave   ctrl
);



endmodule